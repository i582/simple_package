module simple_package

pub fn simple_package_func() int {
    return 0
}
